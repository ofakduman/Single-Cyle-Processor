module xor32(xored, a, b);
	input [31:0]a, b;
	output [31:0]xored;

	xor xoring0(xored[0], a[0], b[0]);
	xor xoring1(xored[1], a[1], b[1]);
	xor xoring2(xored[2], a[2], b[2]);
	xor xoring3(xored[3], a[3], b[3]);
	xor xoring4(xored[4], a[4], b[4]);
	xor xoring5(xored[5], a[5], b[5]);
	xor xoring6(xored[6], a[6], b[6]);
	xor xoring7(xored[7], a[7], b[7]);
	xor xoring8(xored[8], a[8], b[8]);
	xor xoring9(xored[9], a[9], b[9]);
	xor xoring10(xored[10], a[10], b[10]);
	xor xoring11(xored[11], a[11], b[11]);
	xor xoring12(xored[12], a[12], b[12]);
	xor xoring13(xored[13], a[13], b[13]);
	xor xoring14(xored[14], a[14], b[14]);
	xor xoring15(xored[15], a[15], b[15]);
	xor xoring16(xored[16], a[16], b[16]);
	xor xoring17(xored[17], a[17], b[17]);
	xor xoring18(xored[18], a[18], b[18]);
	xor xoring19(xored[19], a[19], b[19]);
	xor xoring20(xored[20], a[20], b[20]);
	xor xoring21(xored[21], a[21], b[21]);
	xor xoring22(xored[22], a[22], b[22]);
	xor xoring23(xored[23], a[23], b[23]);
	xor xoring24(xored[24], a[24], b[24]);
	xor xoring25(xored[25], a[25], b[25]);
	xor xoring26(xored[26], a[26], b[26]);
	xor xoring27(xored[27], a[27], b[27]);
	xor xoring28(xored[28], a[28], b[28]);
	xor xoring29(xored[29], a[29], b[29]);
	xor xoring30(xored[30], a[30], b[30]);
	xor xoring31(xored[31], a[31], b[31]);
endmodule 