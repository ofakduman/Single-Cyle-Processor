module mux_2x1_32(y, op1, op0, s);
input [31:0]op1, op0;
input s;
output [31:0]y;

mux_2x1_1 	m0(y[0],op1[0], op0[0],s),
				m1(y[1],op1[1], op0[1],s),
				m2(y[2],op1[2], op0[2],s),
				m3(y[3],op1[3], op0[3],s),
				m4(y[4],op1[4], op0[4],s),
				m5(y[5],op1[5], op0[5],s),
				m6(y[6],op1[6], op0[6],s),
				m7(y[7],op1[7], op0[7],s),
				m8(y[8],op1[8], op0[8],s),
				m9(y[9],op1[9], op0[9],s),
				m10(y[10],op1[10], op0[10],s),
				m11(y[11],op1[11], op0[11],s),
				m12(y[12],op1[12], op0[12],s),
				m13(y[13],op1[13], op0[13],s),
				m14(y[14],op1[14], op0[14],s),
				m15(y[15],op1[15], op0[15],s),
				m16(y[16],op1[16], op0[16],s),
				m17(y[17],op1[17], op0[17],s),
				m18(y[18],op1[18], op0[18],s),
				m19(y[19],op1[19], op0[19],s),
				m20(y[20],op1[20], op0[20],s),
				m21(y[21],op1[21], op0[21],s),
				m22(y[22],op1[22], op0[22],s),
				m23(y[23],op1[23], op0[23],s),
				m24(y[24],op1[24], op0[24],s),
				m25(y[25],op1[25], op0[25],s),
				m26(y[26],op1[26], op0[26],s),
				m27(y[27],op1[27], op0[27],s),
				m28(y[28],op1[28], op0[28],s),
				m29(y[29],op1[29], op0[29],s),
				m30(y[30],op1[30], op0[30],s),
				m31(y[31],op1[31], op0[31],s);

endmodule
