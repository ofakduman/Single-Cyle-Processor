`define DELAY 100
module alu32_tb(); 

reg [31:0] A,B;
reg [2:0] ALUop;
wire [31:0]R;
wire c_out;
wire signal_reg_write, clk;
wire [31:0] read_data_1,read_data_2;
reg [2:0] read_reg_1, read_reg_2, write_reg,write_data;
wire [31:0] res;
wire Zero0, OverFlow;


alu32 alu(ALUop[2], ALUop[1], ALUop[0], A, B, R, Zero0, OverFlow);

 
initial begin
//ADD
A = 32'b0000_0000_0000_0000_0000_0000_0000_0000; B = 32'b0000_0000_0000_0000_0000_0000_0000_0000; ALUop = 3'b000;
#`DELAY;
A = 32'b0011_0011_0011_0011_0011_0011_0011_0011; B = 32'b0011_0011_0011_0011_0011_0011_0011_0011; ALUop = 3'b000;
#`DELAY;
A = 32'b1111_1111_1111_1111_1111_1111_1111_1111; B = 32'b1111_1111_1111_1111_1111_1111_1111_1111; ALUop = 3'b000;
#`DELAY;
A = 32'b0011_0011_0011_0011_0011_0011_0011_0011; B = 32'b0011_0011_0011_0011_0011_0011_0011_0011; ALUop = 3'b000;
#`DELAY;


//XOR
A = 32'b1000_0001_0001_0010_0010_0101_0000_0000; B = 32'b0000_0000_01110_0000_0000_0000_0000_0000;  ALUop = 3'b001;
#`DELAY;
A = 32'b1011_0011_0011_0011_0011_0011_0011_0011; B = 32'b0011_0011_0011_0011_0011_0011_0011_0011;  ALUop = 3'b001;
#`DELAY;
A = 32'b1011_1011_1111_1001_1101_0011_1111_1011; B = 32'b1111_0001_1111_1111_0000_1111_0011_0011;  ALUop = 3'b001;
#`DELAY;
A = 32'b1010_1111_0011_0001_1011_0010_0000_0011; B = 32'b0011_0011_0011_0011_0011_0111_0011_0011;  ALUop = 3'b001;
#`DELAY;


//SUB
A = 32'b0101_0101_0101_0101_0101_0101_0101_0101; B = 32'b0001_1101_0101_0101_0001_1101_0101_0101;  ALUop = 3'b010;
#`DELAY;
A = 32'b0000_0000_0000_0000_0000_0011_0011_0011; B = 32'b0011_0011_0011_0011_0011_0011_0011_0011;  ALUop = 3'b010;
#`DELAY;
A = 32'b0101_0101_0101_0101_0101_0101_0101_0101; B = 32'b0101_0101_0101_0101_0101_0101_0101_0101;  ALUop = 3'b010;
#`DELAY;
A = 32'b0000_1111_0011_0001_1011_0010_0000_0011; B = 32'b0011_0011_0011_0011_0011_0111_0011_0011;  ALUop = 3'b010;
#`DELAY;


//MULT
A = 32'b1000_0001_0001_0010_0010_0101_0000_0000; B = 32'b0000_0000_0110_0000_0000_0000_0000_0000;  ALUop = 3'b011;
#`DELAY;
A = 32'b1011_0011_0011_0011_0011_0011_0011_0011; B = 32'b0011_0011_0011_0011_0011_0011_0011_0011;  ALUop = 3'b011;
#`DELAY;
A = 32'b1011_1011_1111_1001_1101_0011_1111_1011; B = 32'b1111_0001_1111_1111_0000_1111_0011_0011;  ALUop = 3'b011;
#`DELAY;
A = 32'b1010_1111_0011_0001_1011_0010_0000_0011; B = 32'b0011_0011_0011_0011_0011_0111_0011_0011;  ALUop = 3'b011;
#`DELAY;

//SLT
A = 32'b0101_0101_0101_0101_0101_0101_0101_0101; B = 32'b0001_1101_0101_0101_0001_1101_0101_0101;  ALUop = 3'b100;
#`DELAY;
A = 32'b0000_0000_0000_0000_0000_0011_0011_0011; B = 32'b0011_0011_0011_0011_0011_0011_0011_0011;  ALUop = 3'b100;
#`DELAY;
A = 32'b0101_0101_0101_0101_0101_0101_0101_0101; B = 32'b0101_0101_0101_0101_0101_0101_0101_0101;  ALUop = 3'b100;
#`DELAY;
A = 32'b0000_1111_0011_0001_1011_0010_0000_0011; B = 32'b0011_0011_0011_0011_0011_0111_0011_0011;  ALUop = 3'b100;
#`DELAY;

//NOR
A = 32'b1000_0001_0001_0010_0010_0101_0000_0000; B = 32'b0000_0000_01110_0000_0000_0000_0000_0000;  ALUop = 3'b101;
#`DELAY;
A = 32'b1011_0011_0011_0011_0011_0011_0011_0011; B = 32'b0011_0011_0011_0011_0011_0011_0011_0011;  ALUop = 3'b101;
#`DELAY;
A = 32'b1011_1011_1111_1001_1101_0011_1111_1011; B = 32'b1111_0001_1111_1111_0000_1111_0011_0011;  ALUop = 3'b101;
#`DELAY;
A = 32'b1010_1111_0011_0001_1011_0010_0000_0011; B = 32'b0011_0011_0011_0011_0011_0111_0011_0011;  ALUop = 3'b101;
#`DELAY;


//AND
A = 32'b1000_0001_0001_0010_0010_0101_0000_0000; B = 32'b0000_0000_01110_0000_0000_0000_0000_0000;  ALUop = 3'b110;
#`DELAY;
A = 32'b1011_0011_0011_0011_0011_0011_0011_0011; B = 32'b0011_0011_0011_0011_0011_0011_0011_0011;  ALUop = 3'b110;
#`DELAY;
A = 32'b1011_1011_1111_1001_1101_0011_1111_1011; B = 32'b1111_0001_1111_1111_0000_1111_0011_0011;  ALUop = 3'b110;
#`DELAY;
A = 32'b1010_1111_0011_0001_1011_0010_0000_0011; B = 32'b0011_0011_0011_0011_0011_0111_0011_0011;  ALUop = 3'b110;
#`DELAY;

//OR
A = 32'b1000_0001_0001_0010_0010_0101_0000_0000; B = 32'b0000_0000_01110_0000_0000_0000_0000_0000;  ALUop = 3'b111;
#`DELAY;
A = 32'b1011_0011_0011_0011_0011_0011_0011_0011; B = 32'b0011_0011_0011_0011_0011_0011_0011_0011;  ALUop = 3'b111;
#`DELAY;
A = 32'b1011_1011_1111_1001_1101_0011_1111_1011; B = 32'b1111_0001_1111_1111_0000_1111_0011_0011;  ALUop = 3'b111;
#`DELAY;
A = 32'b1010_1111_0011_0001_1011_0010_0000_0011; B = 32'b0011_0011_0011_0011_0011_0111_0011_0011;  ALUop = 3'b111;
#`DELAY;

end
 
  initial
begin
$monitor("time = %2d, A =%32b, B=%32b, ALUop=%3b, R=%32b",$time, A, B, ALUop, R);
end
 
endmodule